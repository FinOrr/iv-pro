-- Camera registers are reset when there is no power

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity OV5642_Init is
    Port( 
        -- Inputs
        i_Clk       : in  std_logic;
        i_Reset     : in  std_logic;
        i_Next      : in  std_logic;
        -- Outputs
        o_Address   : out  std_logic_vector(15 downto 0);
        o_Data      : out  std_logic_vector(7 downto 0);
        o_Finished  : out  std_logic
    );
end OV5642_Init;

architecture Behavioral of OV5642_Init is
    
    signal r_Reg_Adr : std_logic_vector(15 downto 0) := (x"2FF0");     -- Address of the register we are updating
         
begin
    
    -- Register Reg_Val holds the 8 bit configuration value
    o_Address   <= r_Reg_Adr;
    
    Address_Update: process(i_Clk)
    begin
        if (rising_edge(i_Clk)) then
                if (r_Reg_Adr >= x"589D") then
                    o_Finished <= '1';
                else
                    o_Finished <= '0';
                    if (i_Next = '1') then
                        r_Reg_Adr <= std_logic_vector(unsigned(r_Reg_Adr)+1);
                    end if;
                end if;
            end if;
    end process;
    
    Content_Loader: process(i_Clk)
    begin
        if (rising_edge(i_Clk)) then
            case r_Reg_Adr is
            when x"3000" => o_Data <= x"00";
            when x"3001" => o_Data <= x"00";
            when x"3002" => o_Data <= x"00";
            when x"3003" => o_Data <= x"00";
            when x"3004" => o_Data <= x"ff";
            when x"3008" => o_Data <= x"82";
            when x"300d" => o_Data <= x"22";
            when x"300e" => o_Data <= x"18";
            when x"3010" => o_Data <= x"10";  -- DEF: 00
            when x"3011" => o_Data <= x"08";  -- DEF 14
            when x"3017" => o_Data <= x"7f";
            when x"3018" => o_Data <= x"fc";
            when x"302b" => o_Data <= x"00";
            when x"3030" => o_Data <= x"2b";  -- DEF 0B
            when x"3103" => o_Data <= x"93";
            when x"3406" => o_Data <= x"00";
            when x"3500" => o_Data <= x"00";
            when x"3501" => o_Data <= x"00";
            when x"3502" => o_Data <= x"00";
            when x"3503" => o_Data <= x"00";  -- OR 07
            when x"350a" => o_Data <= x"00";
            when x"350b" => o_Data <= x"00";
            when x"350c" => o_Data <= x"06";
            when x"350d" => o_Data <= x"18";
            when x"3600" => o_Data <= x"52";  -- Analogue control register: 00, 52 or 54
            --when x"3600" => o_Data <= x"54";
            when x"3604" => o_Data <= x"48";
            -- when x"3604" => o_Data <= x"60";
            when x"3605" => o_Data <= x"04";
            -- when x"3606" => o_Data <= x"1b";
            when x"3606" => o_Data <= x"24";
            --  when x"3606" => o_Data <= x"3f";
            when x"3615" => o_Data <= x"f0";
            when x"3620" => o_Data <= x"96";
            when x"3621" => o_Data <= x"10";
            --when x"3621" => o_Data <= x"c9";
            when x"3622" => o_Data <= x"60";
            when x"3623" => o_Data <= x"22";
            when x"3631" => o_Data <= x"01";
            when x"3632" => o_Data <= x"51";
            --   when x"3632" => o_Data <= x"52";
            when x"3702" => o_Data <= x"10";
            when x"3703" => o_Data <= x"b2";
            when x"3704" => o_Data <= x"18";
            when x"3709" => o_Data <= x"00";
            --   when x"3709" => o_Data <= x"01";
            when x"370a" => o_Data <= x"81";
            when x"370b" => o_Data <= x"40";
            when x"370c" => o_Data <= x"a0";
            when x"370d" => o_Data <= x"03";
            when x"370f" => o_Data <= x"c0";
            when x"3710" => o_Data <= x"10";
            when x"3801" => o_Data <= x"88";
            when x"3803" => o_Data <= x"08";
            when x"3804" => o_Data <= x"05";
            when x"3805" => o_Data <= x"00";
            when x"3806" => o_Data <= x"02";
            when x"3807" => o_Data <= x"d0";
            when x"3808" => o_Data <= x"08";  -- or 05
            --when x"3808" => o_Data <= x"0a";
            when x"3809" => o_Data <= x"00";
            when x"380a" => o_Data <= x"06";
            when x"380b" => o_Data <= x"00";
            when x"380c" => o_Data <= x"0c";
            when x"380d" => o_Data <= x"80";
            when x"380e" => o_Data <= x"07";
            when x"380f" => o_Data <= x"d0";
            when x"3810" => o_Data <= x"c2";
            when x"3815" => o_Data <= x"44";
            when x"3818" => o_Data <= x"c9";
            when x"381c" => o_Data <= x"10";
            when x"381d" => o_Data <= x"a0";
            when x"381e" => o_Data <= x"05";
            when x"381f" => o_Data <= x"b0";
            when x"3820" => o_Data <= x"00";
            when x"3821" => o_Data <= x"00";
            when x"3823" => o_Data <= x"00";
            when x"3824" => o_Data <= x"11";
            when x"3825" => o_Data <= x"ac";
            when x"3827" => o_Data <= x"0c";
            when x"3a00" => o_Data <= x"78";
            when x"3a02" => o_Data <= x"00";
            when x"3a03" => o_Data <= x"7d";
            when x"3a04" => o_Data <= x"00";
            when x"3a08" => o_Data <= x"12";
            when x"3a09" => o_Data <= x"c0";
            when x"3a0a" => o_Data <= x"17";
            when x"3a0b" => o_Data <= x"d0";
            when x"3a0d" => o_Data <= x"02";
            when x"3a0e" => o_Data <= x"0d";
            when x"3a0f" => o_Data <= x"30";
            when x"3a10" => o_Data <= x"28";
            when x"3a11" => o_Data <= x"61";
            when x"3a13" => o_Data <= x"30";
            when x"3a14" => o_Data <= x"00";
            when x"3a15" => o_Data <= x"7d";
            when x"3a16" => o_Data <= x"00";
            when x"3a18" => o_Data <= x"00";
            when x"3a19" => o_Data <= x"7c";
            when x"3a1a" => o_Data <= x"04";
            when x"3a1b" => o_Data <= x"30";
            when x"3a1e" => o_Data <= x"28";
            when x"3a1f" => o_Data <= x"10";
            when x"3c00" => o_Data <= x"04";
            when x"3c01" => o_Data <= x"80";
            when x"4000" => o_Data <= x"21";
            when x"4001" => o_Data <= x"42";
            when x"401c" => o_Data <= x"04";
            when x"401d" => o_Data <= x"22";
            when x"401e" => o_Data <= x"20";
            when x"4300" => o_Data <= x"90";
            when x"4402" => o_Data <= x"90";
            when x"4407" => o_Data <= x"04";
            when x"460b" => o_Data <= x"35";
            when x"460c" => o_Data <= x"22";
            when x"4610" => o_Data <= x"00";
            when x"4708" => o_Data <= x"06";
            when x"4713" => o_Data <= x"03";
            when x"471c" => o_Data <= x"50";
            when x"471d" => o_Data <= x"00";
            when x"4721" => o_Data <= x"02";
            when x"5000" => o_Data <= x"df";
            when x"5001" => o_Data <= x"FF";
            when x"5007" => o_Data <= x"00";
            when x"5009" => o_Data <= x"00";
            when x"5011" => o_Data <= x"00";
            when x"5013" => o_Data <= x"00";
            when x"501e" => o_Data <= x"14"; -- Dither ctrl
            when x"501f" => o_Data <= x"00";
            when x"5020" => o_Data <= x"04";
            when x"5025" => o_Data <= x"80";
            when x"5080" => o_Data <= x"08";
            when x"5086" => o_Data <= x"00";
            when x"5087" => o_Data <= x"00";
            when x"5088" => o_Data <= x"00";
            when x"5089" => o_Data <= x"00";
            when x"5180" => o_Data <= x"ff";
            when x"5181" => o_Data <= x"58";
            when x"5182" => o_Data <= x"11";
            when x"5183" => o_Data <= x"14";
            when x"5184" => o_Data <= x"25";
            when x"5185" => o_Data <= x"24";
            when x"5186" => o_Data <= x"14";
            when x"5187" => o_Data <= x"14";
            when x"5188" => o_Data <= x"14";
            when x"5189" => o_Data <= x"69";
            when x"518a" => o_Data <= x"60";
            when x"518b" => o_Data <= x"a2";
            when x"518c" => o_Data <= x"9c";
            when x"518d" => o_Data <= x"36";
            when x"518e" => o_Data <= x"34";
            when x"518f" => o_Data <= x"54";
            when x"5190" => o_Data <= x"4c";
            when x"5191" => o_Data <= x"f8";
            when x"5192" => o_Data <= x"04";
            when x"5193" => o_Data <= x"70";
            when x"5194" => o_Data <= x"f0";
            when x"5195" => o_Data <= x"f0";
            when x"5196" => o_Data <= x"03";
            when x"5197" => o_Data <= x"04";
            when x"5198" => o_Data <= x"05";
            when x"5199" => o_Data <= x"2f";
            when x"519a" => o_Data <= x"04";
            when x"519b" => o_Data <= x"00";
            when x"519c" => o_Data <= x"06";
            when x"519d" => o_Data <= x"a0";
            when x"519e" => o_Data <= x"00";
            when x"5282" => o_Data <= x"00";
            when x"528a" => o_Data <= x"00";
            when x"528b" => o_Data <= x"01";
            when x"528c" => o_Data <= x"04";
            when x"528d" => o_Data <= x"08";
            when x"528e" => o_Data <= x"10";
            when x"528f" => o_Data <= x"20";
            when x"5290" => o_Data <= x"30";
            when x"5292" => o_Data <= x"00";
            when x"5293" => o_Data <= x"00";
            when x"5294" => o_Data <= x"00";
            when x"5295" => o_Data <= x"01";
            when x"5296" => o_Data <= x"00";
            when x"5297" => o_Data <= x"04";
            when x"5298" => o_Data <= x"00";
            when x"5299" => o_Data <= x"08";
            when x"529a" => o_Data <= x"00";
            when x"529b" => o_Data <= x"10";
            when x"529c" => o_Data <= x"00";
            when x"529d" => o_Data <= x"20";
            when x"529e" => o_Data <= x"00";
            when x"529f" => o_Data <= x"30";
            when x"5300" => o_Data <= x"00";
            when x"5301" => o_Data <= x"20";
            when x"5302" => o_Data <= x"00";
            when x"5303" => o_Data <= x"7c";
            when x"5304" => o_Data <= x"00";
            when x"5305" => o_Data <= x"30";
            when x"5306" => o_Data <= x"00";
            when x"5307" => o_Data <= x"80";
            when x"5308" => o_Data <= x"20";
            when x"5309" => o_Data <= x"40";
            when x"530c" => o_Data <= x"00";
            when x"530d" => o_Data <= x"10";
            when x"530e" => o_Data <= x"20";
            when x"530f" => o_Data <= x"80";
            when x"5310" => o_Data <= x"20";
            when x"5311" => o_Data <= x"80";
            when x"5314" => o_Data <= x"08";
            when x"5315" => o_Data <= x"20";
            when x"5316" => o_Data <= x"10";
            when x"5317" => o_Data <= x"00";
            when x"5318" => o_Data <= x"02";
            when x"5319" => o_Data <= x"30";
            when x"5380" => o_Data <= x"01";
            when x"5381" => o_Data <= x"00";
            when x"5382" => o_Data <= x"00";
            when x"5383" => o_Data <= x"1f";
            when x"5384" => o_Data <= x"00";
            when x"5385" => o_Data <= x"06";
            when x"5386" => o_Data <= x"00";
            when x"5387" => o_Data <= x"00";
            when x"5388" => o_Data <= x"00";
            when x"5389" => o_Data <= x"E1";
            when x"538A" => o_Data <= x"00";
            when x"538B" => o_Data <= x"2B";
            when x"538C" => o_Data <= x"00";
            when x"538D" => o_Data <= x"00";
            when x"538E" => o_Data <= x"00";
            when x"538F" => o_Data <= x"10";
            when x"5390" => o_Data <= x"00";
            when x"5391" => o_Data <= x"B3";
            when x"5392" => o_Data <= x"00";
            when x"5393" => o_Data <= x"A6";
            when x"5394" => o_Data <= x"08";
            when x"5402" => o_Data <= x"3f";
            when x"5403" => o_Data <= x"00";
            when x"5480" => o_Data <= x"0c";
            when x"5481" => o_Data <= x"18";
            when x"5482" => o_Data <= x"2f";
            when x"5483" => o_Data <= x"55";
            when x"5484" => o_Data <= x"64";
            when x"5485" => o_Data <= x"71";
            when x"5486" => o_Data <= x"7d";
            when x"5487" => o_Data <= x"87";
            when x"5488" => o_Data <= x"91";
            when x"5489" => o_Data <= x"9a";
            when x"548A" => o_Data <= x"aa";
            when x"548B" => o_Data <= x"b8";
            when x"548C" => o_Data <= x"cd";
            when x"548D" => o_Data <= x"dd";
            when x"548E" => o_Data <= x"ea";
            when x"548F" => o_Data <= x"1d";
            when x"5490" => o_Data <= x"05";
            when x"5491" => o_Data <= x"00";
            when x"5492" => o_Data <= x"04";
            when x"5493" => o_Data <= x"20";
            when x"5494" => o_Data <= x"03";
            when x"5495" => o_Data <= x"60";
            when x"5496" => o_Data <= x"02";
            when x"5497" => o_Data <= x"B8";
            when x"5498" => o_Data <= x"02";
            when x"5499" => o_Data <= x"86";
            when x"549A" => o_Data <= x"02";
            when x"549B" => o_Data <= x"5B";
            when x"549C" => o_Data <= x"02";
            when x"549D" => o_Data <= x"3B";
            when x"549E" => o_Data <= x"02";
            when x"549F" => o_Data <= x"1C";
            when x"54A0" => o_Data <= x"02";
            when x"54A1" => o_Data <= x"04";
            when x"54A2" => o_Data <= x"01";
            when x"54A3" => o_Data <= x"ED";
            when x"54A4" => o_Data <= x"01";
            when x"54A5" => o_Data <= x"C5";
            when x"54A6" => o_Data <= x"01";
            when x"54A7" => o_Data <= x"A5";
            when x"54A8" => o_Data <= x"01";
            when x"54A9" => o_Data <= x"6C";
            when x"54AA" => o_Data <= x"01";
            when x"54AB" => o_Data <= x"41";
            when x"54AC" => o_Data <= x"01";
            when x"54AD" => o_Data <= x"20";
            when x"54AE" => o_Data <= x"00";
            when x"54AF" => o_Data <= x"16";
            when x"54B0" => o_Data <= x"01";
            when x"54B1" => o_Data <= x"20";
            when x"54B2" => o_Data <= x"00";
            when x"54B3" => o_Data <= x"10";
            when x"54B4" => o_Data <= x"00";
            when x"54B5" => o_Data <= x"f0";
            when x"54B6" => o_Data <= x"00";
            when x"54B7" => o_Data <= x"df";
            when x"5500" => o_Data <= x"00";
            when x"5502" => o_Data <= x"00";
            when x"5503" => o_Data <= x"06";
            when x"5504" => o_Data <= x"00";
            when x"5505" => o_Data <= x"FF";
            when x"5580" => o_Data <= x"00";
            when x"5583" => o_Data <= x"40";
            when x"5584" => o_Data <= x"40";
            when x"5682" => o_Data <= x"05";
            when x"5683" => o_Data <= x"00";
            when x"5686" => o_Data <= x"02";
            when x"5687" => o_Data <= x"cc";
            when x"5688" => o_Data <= x"fd";
            when x"5689" => o_Data <= x"df";
            when x"568a" => o_Data <= x"fe";
            when x"568b" => o_Data <= x"ef";
            when x"568c" => o_Data <= x"fe";
            when x"568d" => o_Data <= x"ef";
            when x"568e" => o_Data <= x"aa";
            when x"568f" => o_Data <= x"aa";
            when x"5785" => o_Data <= x"07";
            when x"5800" => o_Data <= x"48";
            when x"5801" => o_Data <= x"31";
            when x"5802" => o_Data <= x"21";
            when x"5803" => o_Data <= x"1b";
            when x"5804" => o_Data <= x"1a";
            when x"5805" => o_Data <= x"1e";
            when x"5806" => o_Data <= x"29";
            when x"5807" => o_Data <= x"38";
            when x"5808" => o_Data <= x"26";
            when x"5809" => o_Data <= x"17";
            when x"580a" => o_Data <= x"11";
            when x"580b" => o_Data <= x"0e";
            when x"580c" => o_Data <= x"0d";
            when x"580d" => o_Data <= x"0e";
            when x"580e" => o_Data <= x"13";
            when x"580f" => o_Data <= x"1a";
            when x"5810" => o_Data <= x"15";
            when x"5811" => o_Data <= x"0d";
            when x"5812" => o_Data <= x"08";
            when x"5813" => o_Data <= x"05";
            when x"5814" => o_Data <= x"04";
            when x"5815" => o_Data <= x"05";
            when x"5816" => o_Data <= x"09";
            when x"5817" => o_Data <= x"0d";
            when x"5818" => o_Data <= x"11";
            when x"5819" => o_Data <= x"0a";
            when x"581a" => o_Data <= x"04";
            when x"581b" => o_Data <= x"00";
            when x"581c" => o_Data <= x"00";
            when x"581d" => o_Data <= x"01";
            when x"581e" => o_Data <= x"06";
            when x"581f" => o_Data <= x"09";
            when x"5820" => o_Data <= x"12";
            when x"5821" => o_Data <= x"0b";
            when x"5822" => o_Data <= x"04";
            when x"5823" => o_Data <= x"00";
            when x"5824" => o_Data <= x"00";
            when x"5825" => o_Data <= x"01";
            when x"5826" => o_Data <= x"06";
            when x"5827" => o_Data <= x"0a";
            when x"5828" => o_Data <= x"17";
            when x"5829" => o_Data <= x"0f";
            when x"582a" => o_Data <= x"09";
            when x"582b" => o_Data <= x"06";
            when x"582c" => o_Data <= x"05";
            when x"582d" => o_Data <= x"06";
            when x"582e" => o_Data <= x"0a";
            when x"582f" => o_Data <= x"0e";
            when x"5830" => o_Data <= x"28";
            when x"5831" => o_Data <= x"1a";
            when x"5832" => o_Data <= x"11";
            when x"5833" => o_Data <= x"0e";
            when x"5834" => o_Data <= x"0e";
            when x"5835" => o_Data <= x"0f";
            when x"5836" => o_Data <= x"15";
            when x"5837" => o_Data <= x"1d";
            when x"5838" => o_Data <= x"6e";
            when x"5839" => o_Data <= x"39";
            when x"583a" => o_Data <= x"27";
            when x"583b" => o_Data <= x"1f";
            when x"583c" => o_Data <= x"1e";
            when x"583d" => o_Data <= x"23";
            when x"583e" => o_Data <= x"2f";
            when x"583f" => o_Data <= x"41";
            when x"5840" => o_Data <= x"0e";
            when x"5841" => o_Data <= x"0c";
            when x"5842" => o_Data <= x"0d";
            when x"5843" => o_Data <= x"0c";
            when x"5844" => o_Data <= x"0c";
            when x"5845" => o_Data <= x"0c";
            when x"5846" => o_Data <= x"0c";
            when x"5847" => o_Data <= x"0c";
            when x"5848" => o_Data <= x"0d";
            when x"5849" => o_Data <= x"0e";
            when x"584a" => o_Data <= x"0e";
            when x"584b" => o_Data <= x"0a";
            when x"584c" => o_Data <= x"0e";
            when x"584d" => o_Data <= x"0e";
            when x"584e" => o_Data <= x"10";
            when x"584f" => o_Data <= x"10";
            when x"5850" => o_Data <= x"11";
            when x"5851" => o_Data <= x"0a";
            when x"5852" => o_Data <= x"0f";
            when x"5853" => o_Data <= x"0e";
            when x"5854" => o_Data <= x"10";
            when x"5855" => o_Data <= x"10";
            when x"5856" => o_Data <= x"10";
            when x"5857" => o_Data <= x"0a";
            when x"5858" => o_Data <= x"0e";
            when x"5859" => o_Data <= x"0e";
            when x"585a" => o_Data <= x"0f";
            when x"585b" => o_Data <= x"0f";
            when x"585c" => o_Data <= x"0f";
            when x"585d" => o_Data <= x"0a";
            when x"585e" => o_Data <= x"09";
            when x"585f" => o_Data <= x"0d";
            when x"5860" => o_Data <= x"0c";
            when x"5861" => o_Data <= x"0b";
            when x"5862" => o_Data <= x"0d";
            when x"5863" => o_Data <= x"07";
            when x"5864" => o_Data <= x"17";
            when x"5865" => o_Data <= x"14";
            when x"5866" => o_Data <= x"18";
            when x"5867" => o_Data <= x"18";
            when x"5868" => o_Data <= x"16";
            when x"5869" => o_Data <= x"12";
            when x"586a" => o_Data <= x"1b";
            when x"586b" => o_Data <= x"1a";
            when x"586c" => o_Data <= x"16";
            when x"586d" => o_Data <= x"16";
            when x"586e" => o_Data <= x"18";
            when x"586f" => o_Data <= x"1f";
            when x"5870" => o_Data <= x"1c";
            when x"5871" => o_Data <= x"16";
            when x"5872" => o_Data <= x"10";
            when x"5873" => o_Data <= x"0f";
            when x"5874" => o_Data <= x"13";
            when x"5875" => o_Data <= x"1c";
            when x"5876" => o_Data <= x"1e";
            when x"5877" => o_Data <= x"17";
            when x"5878" => o_Data <= x"11";
            when x"5879" => o_Data <= x"11";
            when x"587a" => o_Data <= x"14";
            when x"587b" => o_Data <= x"1e";
            when x"587c" => o_Data <= x"1c";
            when x"587d" => o_Data <= x"1c";
            when x"587e" => o_Data <= x"1a";
            when x"587f" => o_Data <= x"1a";
            when x"5880" => o_Data <= x"1b";
            when x"5881" => o_Data <= x"1f";
            when x"5882" => o_Data <= x"14";
            when x"5883" => o_Data <= x"1a";
            when x"5884" => o_Data <= x"1d";
            when x"5885" => o_Data <= x"1e";
            when x"5886" => o_Data <= x"1a";
            when x"5887" => o_Data <= x"1a";
            when x"589a" => o_Data <= x"c0";
            when x"589b" => o_Data <= x"00";
            when others  => o_Data <= (others => 'Z');
            end case;
        end if;
    end process;
end Behavioral;